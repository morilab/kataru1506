/////////////////////////////////////////////////////////////////////////////
// Engineer      : $Author: MoriLab. $
// Create Date   : 2013/03/30 12:00:00
// Design Name   : $RCSfile: packet.svh,v $
// Project Name  : Packet
// Project No.   : 
// Syntax        : OVM2.0.3
// Tool versions : ModelSim10.1
// Revision      : $Revision: 1.1 $
// Last Update   : $Date: 2013/04/11 00:35:11 $ + 09:00:00
//<Additional Comments>//////////////////////////////////////////////////////
///
/////////////////////////////////////////////////////////////////////////////
package ovm_Packet_pkg;
	`include "vt100.svh"
	`include "ovm_macros.svh"
	import ovm_pkg::*;
	`include "packet_item.sv"
endpackage
