/////////////////////////////////////////////////////////////////////////////
// Engineer      : $Author: MoriLab. $
// Create Date   : Wed, 17 Jun 2015 01:47:38 +0900 
// Design Name   : $RCSfile: verienv_apb2iic_test_list.sv,v $
// Project Name  : kataru1506 
// Project No.   : - 
// Syntax        : ovm-2.0.3
// Tool versions : Model Technology ModelSim ALTERA STARTER EDITION vsim 10.1d Simulator 2012.11 Nov 2 2012
// Revision      : $Revision: 1.3 $
// Last Update   : $Date: 2012/03/26 12:20:12 $ + 09:00:00
//<Additional Comments>//////////////////////////////////////////////////////
// �e�X�g���ꗗ
/////////////////////////////////////////////////////////////////////////////

// �e�X�g��
`include "test/verienv_apb2iic_test0001_test.sv"
`include "test/verienv_apb2iic_test0002_test.sv"
//TEST//

// �e�X�g�V�i���I
`include "test/verienv_apb2iic_test0001_vseq.sv"
`include "test/verienv_apb2iic_test0002_vseq.sv"
//VSEQ//

