/////////////////////////////////////////////////////////////////////////////
// Engineer      : $Author: MoriLab. $
// Create Date   : Wed, 17 Jun 2015 01:47:38 +0900 
// Design Name   : $RCSfile: tb_top.sv,v $
// Project Name  : kataru1506 
// Project No.   : - 
// Syntax        : ovm-2.0.3
// Tool versions : Model Technology ModelSim ALTERA STARTER EDITION vsim 10.1d Simulator 2012.11 Nov 2 2012
// Revision      : $Revision: 1.3 $
// Last Update   : $Date: 2012/10/19 13:13:44 $ + 09:00:00
//<Additional Comments>//////////////////////////////////////////////////////
// ���؊����W���[��
// �S�̌��؊�
/////////////////////////////////////////////////////////////////////////////
// OVM�W�����C�u����

// �C���^�[�t�F�[�X�錾

// ���b�p�[
/// ���؃g�b�v���W���[��
module tb_top();
	
	// OVM���f�����C�u����
	
	// �^�錾
	
	// �C���^�[�t�F�[�X
	
	// ����RTL�g�b�v
	DUV DUV (                                 // <DUV>
	);                                        // </>
endmodule
