/////////////////////////////////////////////////////////////////////////////
// Engineer      : $Author: MoriLab. $
// Create Date   : Wed, 17 Jun 2015 01:47:38 +0900 
// Design Name   : $RCSfile: tb_top.sv,v $
// Project Name  : kataru1506 
// Project No.   : - 
// Syntax        : ovm-2.0.3
// Tool versions : Model Technology ModelSim ALTERA STARTER EDITION vsim 10.1d Simulator 2012.11 Nov 2 2012
// Revision      : $Revision: 1.3 $
// Last Update   : $Date: 2012/10/19 13:13:44 $ + 09:00:00
//<Additional Comments>//////////////////////////////////////////////////////
// 検証環境モジュール
// 全体検証環境
/////////////////////////////////////////////////////////////////////////////
// OVM標準ライブラリ

// インターフェース宣言

// ラッパー
/// 検証トップモジュール
module tb_top();
	
	// OVMモデルライブラリ
	
	// 型宣言
	
	// インターフェース
	
	// 検証RTLトップ
	DUV DUV (                                 // <DUV>
	);                                        // </>
endmodule
