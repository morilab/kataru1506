/////////////////////////////////////////////////////////////////////////////
// Engineer      : $Author: MoriLab. $
// Create Date   : 2012/01/19 12:00:00
// Design Name   : $RCSfile: scoreboard_share.sv,v $
// Project Name  : ScoreBoard
// Project No.   : 
// Syntax        : OVM2.0.3
// Tool versions : ModelSim10.1
// Revision      : $Revision: 1.1 $
// Last Update   : $Date: 2012/03/26 05:38:31 $ + 09:00:00
//<Additional Comments>//////////////////////////////////////////////////////
// ��ͭ�ѿ�
/////////////////////////////////////////////////////////////////////////////

///@brief   �����å��⡼��
///@details �������ܡ��ɤǼ������������ƥ�Υ����å���ˡ�򼨤��ޤ���
typedef enum {
	IN_ORDER   , ///< ���󥪡��������
	OUT_ORDER  , ///< �����ȥ����������
	COUNT_ONLY , ///< ���Τߤ����
	NO_COMPARE   ///< ��Ӥ��ʤ�
} chk_rule;

///@brief   �������
///@details ��������η��򼨤��ޤ���
///@warning ���ε�ǽ�Ͼ���Ū�˼�������٤��Ǥ��������ߤ�̤�����Ǥ���
///@note    ưŪ����ϥ��������Ϲ�®�Ǥ��������ɥ쥹������ʬ�Υ������ݤ����1MB��Ķ����褦�ʶ��֤ˤϸ����ޤ���
///         Ϣ������ϥ���������ưŪ�������٤����®�Ǥ��������������������ɥ쥹�˴ؤ��ƤΤߡʥ����������������ǡ�
///         �������ݤ���١��������ɥ쥹���֤ΰ����Τߥ�����������褦��ư���Ŭ���Ƥ��ޤ���<br>
///         �����ߤ�Ϣ������ˤ�������ԤäƤ��ޤ���
typedef enum {
	RAM_IS_DYNAMIC_ARRAY     , ///< ưŪ����
	RAM_IS_ASSOCIATIVE_ARRAY   ///< Ϣ������
} sb_ram_type;
